class spi_transaction extend uvm_sequence_item;


endclass