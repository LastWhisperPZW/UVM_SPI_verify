it remote add origin git@github.com:LastWhisperPZW/UVM_SPI_verify
