`ifndef SPI_TRANSACTION__SV
`define SPI_TRANSACTION__SV

class spi_transaction extends uvm_sequence_item;


endclass

`endif