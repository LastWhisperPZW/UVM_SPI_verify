uvm_env extends